module mips_ex (
);



endmodule // EXU
